module vmujs

fn test_simple_function() {
	assert false
}
